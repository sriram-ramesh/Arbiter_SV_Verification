//                              -*- Mode: Verilog -*-
// Filename        : scoreboard.sv
// Description     : scoreboard for arbiter
// Author          : vinchip
// Created On      : Mon Aug 24 17:34:27 2015
// Last Modified By: .
// Last Modified On: .
// Update Count    : 0
// Status          : Unknown, Use with caution!
/////////////////////////////////////////////////////


class scoreboard;
   
   bit grant1,grant2,grant3,grant4;
   
   

endclass // scoreboard
